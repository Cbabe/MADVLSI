magic
tech sky130A
timestamp 1695933658
<< nwell >>
rect -315 315 -225 435
rect -45 315 180 580
rect -575 165 180 315
rect -575 10 -365 165
rect -575 5 -380 10
<< nmos >>
rect -145 490 -130 590
rect -145 360 -130 460
rect -315 -130 -300 -30
rect -245 -130 -230 -30
rect 25 -130 40 -30
rect 95 -130 110 -30
rect -315 -385 -300 -185
<< pmos >>
rect 75 355 90 555
rect -470 155 -455 255
rect -315 185 -300 285
rect -245 185 -230 285
rect 25 185 40 285
rect 95 185 110 285
rect -470 25 -455 125
<< ndiff >>
rect -190 575 -145 590
rect -190 505 -180 575
rect -160 505 -145 575
rect -190 490 -145 505
rect -130 575 -80 590
rect -130 505 -115 575
rect -95 505 -80 575
rect -130 490 -80 505
rect -190 445 -145 460
rect -190 375 -180 445
rect -160 375 -145 445
rect -190 360 -145 375
rect -130 445 -80 460
rect -130 375 -115 445
rect -95 375 -80 445
rect -130 360 -80 375
rect -365 -45 -315 -30
rect -365 -115 -350 -45
rect -330 -115 -315 -45
rect -365 -130 -315 -115
rect -300 -45 -245 -30
rect -300 -115 -285 -45
rect -265 -115 -245 -45
rect -300 -130 -245 -115
rect -230 -45 -180 -30
rect -230 -115 -215 -45
rect -195 -115 -180 -45
rect -230 -130 -180 -115
rect -25 -45 25 -30
rect -25 -115 -10 -45
rect 10 -115 25 -45
rect -25 -130 25 -115
rect 40 -45 95 -30
rect 40 -115 55 -45
rect 75 -115 95 -45
rect 40 -130 95 -115
rect 110 -45 160 -30
rect 110 -115 125 -45
rect 145 -115 160 -45
rect 110 -130 160 -115
rect -365 -200 -315 -185
rect -365 -370 -350 -200
rect -330 -370 -315 -200
rect -365 -385 -315 -370
rect -300 -200 -245 -185
rect -300 -370 -285 -200
rect -265 -370 -245 -200
rect -300 -385 -245 -370
<< pdiff >>
rect 30 540 75 555
rect 30 370 40 540
rect 60 370 75 540
rect 30 355 75 370
rect 90 540 140 555
rect 90 370 105 540
rect 125 370 140 540
rect 90 355 140 370
rect -365 270 -315 285
rect -515 240 -470 255
rect -515 170 -505 240
rect -485 170 -470 240
rect -515 155 -470 170
rect -455 240 -405 255
rect -455 170 -440 240
rect -420 170 -405 240
rect -365 200 -350 270
rect -330 200 -315 270
rect -365 185 -315 200
rect -300 270 -245 285
rect -300 200 -285 270
rect -265 200 -245 270
rect -300 185 -245 200
rect -230 270 -180 285
rect -230 200 -215 270
rect -195 200 -180 270
rect -230 185 -180 200
rect -25 270 25 285
rect -25 200 -10 270
rect 10 200 25 270
rect -25 185 25 200
rect 40 270 95 285
rect 40 200 55 270
rect 75 200 95 270
rect 40 185 95 200
rect 110 270 160 285
rect 110 200 125 270
rect 145 200 160 270
rect 110 185 160 200
rect -455 155 -405 170
rect -515 110 -470 125
rect -515 40 -505 110
rect -485 40 -470 110
rect -515 25 -470 40
rect -455 110 -405 125
rect -455 40 -440 110
rect -420 40 -405 110
rect -455 25 -405 40
<< ndiffc >>
rect -180 505 -160 575
rect -115 505 -95 575
rect -180 375 -160 445
rect -115 375 -95 445
rect -350 -115 -330 -45
rect -285 -115 -265 -45
rect -215 -115 -195 -45
rect -10 -115 10 -45
rect 55 -115 75 -45
rect 125 -115 145 -45
rect -350 -370 -330 -200
rect -285 -370 -265 -200
<< pdiffc >>
rect 40 370 60 540
rect 105 370 125 540
rect -505 170 -485 240
rect -440 170 -420 240
rect -350 200 -330 270
rect -285 200 -265 270
rect -215 200 -195 270
rect -10 200 10 270
rect 55 200 75 270
rect 125 200 145 270
rect -505 40 -485 110
rect -440 40 -420 110
<< psubdiff >>
rect 45 -175 95 -160
rect -415 -200 -365 -185
rect -415 -370 -400 -200
rect -380 -370 -365 -200
rect -415 -385 -365 -370
rect 45 -245 60 -175
rect 80 -245 95 -175
rect 45 -260 95 -245
<< nsubdiff >>
rect -20 540 30 555
rect -295 400 -245 415
rect -295 330 -280 400
rect -260 330 -245 400
rect -20 370 -5 540
rect 15 370 30 540
rect -20 355 30 370
rect -295 315 -245 330
<< psubdiffcont >>
rect -400 -370 -380 -200
rect 60 -245 80 -175
<< nsubdiffcont >>
rect -280 330 -260 400
rect -5 370 15 540
<< poly >>
rect -575 600 180 615
rect -470 255 -455 600
rect -145 590 -130 600
rect 75 555 90 600
rect -145 460 -130 490
rect -145 345 -130 360
rect 75 340 90 355
rect -125 315 -85 320
rect -125 310 40 315
rect -315 285 -300 300
rect -245 285 -230 300
rect -125 290 -115 310
rect -95 300 40 310
rect -95 290 -85 300
rect -125 280 -85 290
rect 25 285 40 300
rect 95 285 110 300
rect -470 125 -455 155
rect -380 120 -340 130
rect -380 100 -370 120
rect -350 100 -340 120
rect -380 90 -340 100
rect -375 30 -360 90
rect -315 70 -300 185
rect -245 135 -230 185
rect -270 125 -230 135
rect -205 160 -165 170
rect -205 140 -195 160
rect -175 140 -165 160
rect -205 130 -165 140
rect -270 105 -260 125
rect -240 105 -230 125
rect -270 95 -230 105
rect -315 60 -275 70
rect -315 40 -305 60
rect -285 40 -275 60
rect -315 30 -275 40
rect -470 -395 -455 25
rect -380 20 -340 30
rect -380 0 -370 20
rect -350 0 -340 20
rect -380 -10 -340 0
rect -315 -30 -300 30
rect -245 -30 -230 95
rect -190 70 -175 130
rect -40 120 0 130
rect -40 100 -30 120
rect -10 100 0 120
rect -40 90 0 100
rect -205 60 -165 70
rect -205 40 -195 60
rect -175 40 -165 60
rect -205 30 -165 40
rect -35 30 -20 90
rect 25 70 40 185
rect 95 135 110 185
rect 70 125 110 135
rect 135 160 175 170
rect 135 140 145 160
rect 165 140 175 160
rect 135 130 175 140
rect 70 105 80 125
rect 100 105 110 125
rect 70 95 110 105
rect 25 60 65 70
rect 25 40 35 60
rect 55 40 65 60
rect 25 30 65 40
rect -40 20 0 30
rect -40 0 -30 20
rect -10 0 0 20
rect -40 -10 0 0
rect 25 -30 40 30
rect 95 -30 110 95
rect 150 70 165 130
rect 135 60 175 70
rect 135 40 145 60
rect 165 40 175 60
rect 135 30 175 40
rect -315 -145 -300 -130
rect -245 -145 -230 -130
rect 25 -145 40 -130
rect 95 -145 110 -130
rect -315 -185 -300 -170
rect -315 -395 -300 -385
rect -470 -410 -300 -395
<< polycont >>
rect -115 290 -95 310
rect -370 100 -350 120
rect -195 140 -175 160
rect -260 105 -240 125
rect -305 40 -285 60
rect -370 0 -350 20
rect -30 100 -10 120
rect -195 40 -175 60
rect 145 140 165 160
rect 80 105 100 125
rect 35 40 55 60
rect -30 0 -10 20
rect 145 40 165 60
<< locali >>
rect -190 575 -150 585
rect -190 515 -180 575
rect -340 505 -180 515
rect -160 505 -150 575
rect -340 495 -150 505
rect -125 575 -85 585
rect -125 505 -115 575
rect -95 515 -85 575
rect -20 540 70 550
rect -95 505 -40 515
rect -125 495 -40 505
rect -340 280 -320 495
rect -190 445 -150 455
rect -290 400 -250 410
rect -290 330 -280 400
rect -260 330 -250 400
rect -190 385 -180 445
rect -290 320 -250 330
rect -205 375 -180 385
rect -160 375 -150 445
rect -205 365 -150 375
rect -125 445 -85 455
rect -125 375 -115 445
rect -95 375 -85 445
rect -125 365 -85 375
rect -275 280 -255 320
rect -205 280 -185 365
rect -115 320 -95 365
rect -60 340 -40 495
rect -20 370 -5 540
rect 15 370 40 540
rect 60 370 70 540
rect -20 360 70 370
rect 95 540 135 550
rect 95 370 105 540
rect 125 370 135 540
rect 95 360 135 370
rect -60 320 -5 340
rect 105 335 125 360
rect 70 325 125 335
rect -125 310 -85 320
rect -125 290 -115 310
rect -95 290 -85 310
rect -125 280 -85 290
rect -25 280 -5 320
rect 65 315 125 325
rect 65 280 85 315
rect -365 270 -320 280
rect -515 240 -475 250
rect -515 180 -505 240
rect -555 170 -505 180
rect -485 170 -475 240
rect -555 160 -475 170
rect -450 240 -410 250
rect -450 170 -440 240
rect -420 180 -410 240
rect -365 200 -350 270
rect -330 200 -320 270
rect -365 190 -320 200
rect -295 270 -255 280
rect -295 200 -285 270
rect -265 200 -255 270
rect -295 190 -255 200
rect -225 270 -185 280
rect -225 200 -215 270
rect -195 200 -185 270
rect -225 190 -185 200
rect -365 180 -345 190
rect -420 170 -345 180
rect -450 160 -345 170
rect -555 110 -535 160
rect -365 130 -345 160
rect -205 170 -185 190
rect -25 270 20 280
rect -25 200 -10 270
rect 10 200 20 270
rect -25 190 20 200
rect 45 270 85 280
rect 45 200 55 270
rect 75 200 85 270
rect 45 190 85 200
rect 115 270 155 280
rect 115 200 125 270
rect 145 200 155 270
rect 115 190 155 200
rect -205 160 -165 170
rect -205 140 -195 160
rect -175 140 -165 160
rect -380 120 -340 130
rect -270 125 -230 135
rect -205 130 -165 140
rect -25 130 -5 190
rect 135 170 155 190
rect 135 160 175 170
rect 135 140 145 160
rect 165 140 175 160
rect -270 120 -260 125
rect -575 90 -535 110
rect -510 110 -475 120
rect -510 70 -505 110
rect -575 50 -505 70
rect -535 45 -505 50
rect -510 40 -505 45
rect -485 40 -475 110
rect -510 30 -475 40
rect -450 110 -410 120
rect -450 40 -440 110
rect -420 70 -410 110
rect -380 100 -370 120
rect -350 110 -340 120
rect -290 110 -260 120
rect -350 105 -260 110
rect -240 105 -230 125
rect -350 100 -230 105
rect -380 95 -230 100
rect -40 120 0 130
rect 70 125 110 135
rect 135 130 175 140
rect 70 120 80 125
rect -40 100 -30 120
rect -10 110 0 120
rect 50 110 80 120
rect -10 105 80 110
rect 100 120 110 125
rect 100 115 115 120
rect 100 110 125 115
rect 100 105 180 110
rect -10 100 180 105
rect -40 95 180 100
rect -380 90 -280 95
rect -40 90 60 95
rect 110 90 180 95
rect -420 60 -165 70
rect -420 50 -305 60
rect -420 40 -410 50
rect -450 30 -410 40
rect -315 40 -305 50
rect -285 50 -195 60
rect -285 40 -275 50
rect -315 30 -275 40
rect -205 40 -195 50
rect -175 40 -165 60
rect -35 60 180 70
rect -35 50 35 60
rect -205 30 -165 40
rect 25 40 35 50
rect 55 50 145 60
rect 55 40 65 50
rect 25 30 65 40
rect 135 40 145 50
rect 165 45 180 60
rect 165 40 175 45
rect 135 30 175 40
rect -380 20 -340 30
rect -380 0 -370 20
rect -350 0 -340 20
rect -380 -10 -340 0
rect -365 -35 -345 -10
rect -205 -35 -185 30
rect -40 20 0 30
rect -40 0 -30 20
rect -10 0 0 20
rect -40 -10 0 0
rect -365 -45 -320 -35
rect -365 -115 -350 -45
rect -330 -115 -320 -45
rect -365 -125 -320 -115
rect -295 -45 -250 -35
rect -295 -115 -285 -45
rect -265 -115 -250 -45
rect -295 -125 -250 -115
rect -225 -45 -185 -35
rect -225 -115 -215 -45
rect -195 -115 -185 -45
rect -225 -125 -185 -115
rect -25 -35 -5 -10
rect 135 -35 155 30
rect -25 -45 20 -35
rect -25 -115 -10 -45
rect 10 -115 20 -45
rect -25 -125 20 -115
rect 45 -45 90 -35
rect 45 -115 55 -45
rect 75 -115 90 -45
rect 45 -125 90 -115
rect 115 -45 155 -35
rect 115 -115 125 -45
rect 145 -115 155 -45
rect 115 -125 155 -115
rect -280 -190 -260 -125
rect 60 -165 80 -125
rect 45 -175 95 -165
rect -415 -200 -320 -190
rect -415 -370 -400 -200
rect -380 -370 -350 -200
rect -330 -370 -320 -200
rect -415 -380 -320 -370
rect -295 -200 -250 -190
rect -295 -370 -285 -200
rect -265 -370 -250 -200
rect 45 -245 60 -175
rect 80 -245 95 -175
rect 45 -255 95 -245
rect -295 -380 -250 -370
rect -280 -385 -260 -380
<< viali >>
rect -280 330 -260 400
rect -5 370 15 540
rect -400 -370 -380 -200
rect 60 -245 80 -175
<< metal1 >>
rect -190 550 -80 585
rect -575 540 180 550
rect -575 400 -5 540
rect -575 330 -280 400
rect -260 370 -5 400
rect 15 370 180 540
rect -260 330 180 370
rect -575 320 180 330
rect -295 315 -245 320
rect -575 -175 180 -165
rect -575 -200 60 -175
rect -575 -370 -400 -200
rect -380 -245 60 -200
rect 80 -245 180 -175
rect -380 -370 180 -245
rect -575 -400 180 -370
<< labels >>
rlabel metal1 -575 445 -575 445 7 VDD
port 4 w
rlabel metal1 -575 -255 -575 -255 7 GND
port 1 w
rlabel locali -575 60 -575 60 7 D_bar
port 2 w
rlabel locali -575 100 -575 100 7 D
port 3 w
rlabel poly -575 605 -575 605 7 Phi
port 5 w
rlabel locali 180 55 180 55 3 Q_bar
port 7 e
rlabel locali 180 100 180 100 3 Q
port 6 e
<< end >>
