magic
tech sky130A
timestamp 1695938287
<< error_p >>
rect -228 885 -205 903
rect -145 885 -101 969
rect -228 875 -101 885
rect -210 855 -101 875
rect -210 824 -151 855
rect -235 808 -151 824
rect -253 785 -151 808
rect -253 767 -192 785
<< nwell >>
rect -360 1450 -110 1600
rect -360 1255 -135 1450
rect -365 1185 -135 1255
rect -365 1135 -145 1185
rect -370 1125 -145 1135
rect -375 885 -145 1125
rect -375 855 -210 885
rect -185 855 -145 885
rect -235 785 -210 855
rect -315 360 -225 435
rect -375 315 -225 360
rect -375 305 -205 315
rect -375 300 -160 305
rect -385 270 -160 300
rect -400 165 -160 270
<< nmos >>
rect -290 1795 -275 1895
rect -220 1795 -205 1895
rect -270 690 -255 790
rect -270 560 -255 660
rect -315 -130 -300 -30
rect -245 -130 -230 -30
rect -315 -385 -300 -185
<< pmos >>
rect -290 1480 -275 1580
rect -220 1480 -205 1580
rect -270 1210 -255 1410
rect -270 1005 -255 1105
rect -270 875 -255 975
rect -315 185 -300 285
rect -245 185 -230 285
<< ndiff >>
rect -340 1880 -290 1895
rect -340 1810 -325 1880
rect -305 1810 -290 1880
rect -340 1795 -290 1810
rect -275 1880 -220 1895
rect -275 1810 -255 1880
rect -235 1810 -220 1880
rect -275 1795 -220 1810
rect -205 1880 -155 1895
rect -205 1810 -190 1880
rect -170 1810 -155 1880
rect -205 1795 -155 1810
rect -315 775 -270 790
rect -315 705 -305 775
rect -285 705 -270 775
rect -315 690 -270 705
rect -255 785 -235 790
rect -210 785 -205 790
rect -255 775 -205 785
rect -255 705 -240 775
rect -220 705 -205 775
rect -255 690 -205 705
rect -315 645 -270 660
rect -315 585 -305 645
rect -310 575 -305 585
rect -285 575 -270 645
rect -310 560 -270 575
rect -255 645 -205 660
rect -255 575 -240 645
rect -220 575 -205 645
rect -255 560 -205 575
rect -365 -45 -315 -30
rect -365 -115 -350 -45
rect -330 -115 -315 -45
rect -365 -130 -315 -115
rect -300 -45 -245 -30
rect -300 -115 -285 -45
rect -265 -115 -245 -45
rect -300 -130 -245 -115
rect -230 -45 -180 -30
rect -230 -115 -215 -45
rect -195 -115 -180 -45
rect -230 -130 -180 -115
rect -365 -200 -315 -185
rect -365 -370 -350 -200
rect -330 -370 -315 -200
rect -365 -385 -315 -370
rect -300 -200 -245 -185
rect -300 -370 -285 -200
rect -265 -370 -245 -200
rect -300 -385 -245 -370
<< pdiff >>
rect -340 1565 -290 1580
rect -340 1495 -325 1565
rect -305 1495 -290 1565
rect -340 1480 -290 1495
rect -275 1565 -220 1580
rect -275 1495 -255 1565
rect -235 1495 -220 1565
rect -275 1480 -220 1495
rect -205 1565 -155 1580
rect -205 1495 -190 1565
rect -170 1495 -155 1565
rect -205 1480 -155 1495
rect -320 1395 -270 1410
rect -320 1225 -305 1395
rect -285 1225 -270 1395
rect -320 1210 -270 1225
rect -255 1395 -210 1410
rect -255 1225 -240 1395
rect -220 1225 -210 1395
rect -255 1210 -210 1225
rect -315 1090 -270 1105
rect -315 1020 -305 1090
rect -285 1020 -270 1090
rect -315 1005 -270 1020
rect -255 1090 -205 1105
rect -255 1020 -240 1090
rect -220 1020 -205 1090
rect -255 1005 -205 1020
rect -315 960 -270 975
rect -315 890 -305 960
rect -285 890 -270 960
rect -315 875 -270 890
rect -255 960 -205 975
rect -255 890 -240 960
rect -220 890 -205 960
rect -255 885 -205 890
rect -255 875 -210 885
rect -235 785 -210 790
rect -365 270 -315 285
rect -365 200 -350 270
rect -330 200 -315 270
rect -365 185 -315 200
rect -300 270 -245 285
rect -300 200 -285 270
rect -265 200 -245 270
rect -300 185 -245 200
rect -230 270 -180 285
rect -230 200 -215 270
rect -195 200 -180 270
rect -230 185 -180 200
<< ndiffc >>
rect -325 1810 -305 1880
rect -255 1810 -235 1880
rect -190 1810 -170 1880
rect -305 705 -285 775
rect -240 705 -220 775
rect -305 575 -285 645
rect -240 575 -220 645
rect -350 -115 -330 -45
rect -285 -115 -265 -45
rect -215 -115 -195 -45
rect -350 -370 -330 -200
rect -285 -370 -265 -200
<< pdiffc >>
rect -325 1495 -305 1565
rect -255 1495 -235 1565
rect -190 1495 -170 1565
rect -305 1225 -285 1395
rect -240 1225 -220 1395
rect -305 1020 -285 1090
rect -240 1020 -220 1090
rect -305 890 -285 960
rect -240 890 -220 960
rect -350 200 -330 270
rect -285 200 -265 270
rect -215 200 -195 270
<< psubdiff >>
rect -275 2010 -225 2025
rect -275 1940 -260 2010
rect -240 1940 -225 2010
rect -275 1925 -225 1940
rect -415 -200 -365 -185
rect -415 -370 -400 -200
rect -380 -370 -365 -200
rect -415 -385 -365 -370
<< nsubdiff >>
rect -210 1395 -160 1410
rect -210 1225 -195 1395
rect -175 1225 -160 1395
rect -210 1210 -160 1225
rect -295 400 -245 415
rect -295 330 -280 400
rect -260 330 -245 400
rect -295 315 -245 330
<< psubdiffcont >>
rect -260 1940 -240 2010
rect -400 -370 -380 -200
<< nsubdiffcont >>
rect -195 1225 -175 1395
rect -280 330 -260 400
<< poly >>
rect -290 1895 -275 1910
rect -220 1895 -205 1910
rect -355 1725 -315 1735
rect -355 1705 -345 1725
rect -325 1705 -315 1725
rect -355 1695 -315 1705
rect -345 1635 -330 1695
rect -290 1670 -275 1795
rect -220 1735 -205 1795
rect -180 1765 -140 1775
rect -180 1745 -170 1765
rect -150 1745 -140 1765
rect -180 1735 -140 1745
rect -245 1725 -205 1735
rect -245 1705 -235 1725
rect -215 1705 -205 1725
rect -245 1695 -205 1705
rect -290 1660 -250 1670
rect -290 1640 -280 1660
rect -260 1640 -250 1660
rect -355 1625 -315 1635
rect -355 1605 -345 1625
rect -325 1605 -315 1625
rect -355 1595 -315 1605
rect -290 1630 -250 1640
rect -290 1580 -275 1630
rect -220 1580 -205 1695
rect -160 1675 -145 1735
rect -180 1665 -140 1675
rect -180 1645 -170 1665
rect -150 1645 -140 1665
rect -180 1635 -140 1645
rect -290 1465 -275 1480
rect -220 1465 -205 1480
rect -220 1450 -95 1465
rect -270 1410 -255 1425
rect -270 1105 -255 1210
rect -110 1185 -95 1450
rect -270 975 -255 1005
rect -270 790 -255 875
rect -185 815 -180 835
rect -270 660 -255 690
rect -270 545 -255 560
rect -440 530 -255 545
rect -440 -395 -425 530
rect -185 520 -170 815
rect -225 510 -170 520
rect -225 490 -215 510
rect -195 500 -170 510
rect -195 490 -185 500
rect -225 480 -185 490
rect -315 285 -300 300
rect -245 285 -230 300
rect -380 120 -340 130
rect -380 100 -370 120
rect -350 100 -340 120
rect -380 90 -340 100
rect -375 30 -360 90
rect -315 70 -300 185
rect -245 135 -230 185
rect -270 125 -230 135
rect -205 160 -165 170
rect -205 140 -195 160
rect -175 140 -165 160
rect -205 130 -165 140
rect -270 105 -260 125
rect -240 105 -230 125
rect -270 95 -230 105
rect -315 60 -275 70
rect -315 40 -305 60
rect -285 40 -275 60
rect -315 30 -275 40
rect -380 20 -340 30
rect -380 0 -370 20
rect -350 0 -340 20
rect -380 -10 -340 0
rect -315 -30 -300 30
rect -245 -30 -230 95
rect -190 70 -175 130
rect -205 60 -165 70
rect -205 40 -195 60
rect -175 40 -165 60
rect -205 30 -165 40
rect -315 -145 -300 -130
rect -245 -145 -230 -130
rect -315 -185 -300 -170
rect -315 -395 -300 -385
rect -440 -410 -300 -395
<< polycont >>
rect -345 1705 -325 1725
rect -170 1745 -150 1765
rect -235 1705 -215 1725
rect -280 1640 -260 1660
rect -345 1605 -325 1625
rect -170 1645 -150 1665
rect -215 490 -195 510
rect -370 100 -350 120
rect -195 140 -175 160
rect -260 105 -240 125
rect -305 40 -285 60
rect -370 0 -350 20
rect -195 40 -175 60
<< locali >>
rect -275 2010 -225 2020
rect -275 1940 -260 2010
rect -240 1940 -225 2010
rect -275 1930 -225 1940
rect -260 1890 -240 1930
rect -335 1880 -295 1890
rect -335 1810 -325 1880
rect -305 1810 -295 1880
rect -335 1800 -295 1810
rect -270 1880 -225 1890
rect -270 1810 -255 1880
rect -235 1810 -225 1880
rect -270 1800 -225 1810
rect -200 1880 -155 1890
rect -200 1810 -190 1880
rect -170 1810 -155 1880
rect -200 1800 -155 1810
rect -335 1735 -315 1800
rect -175 1775 -155 1800
rect -180 1765 -140 1775
rect -180 1745 -170 1765
rect -150 1745 -140 1765
rect -180 1735 -140 1745
rect -355 1725 -315 1735
rect -355 1720 -345 1725
rect -360 1705 -345 1720
rect -325 1715 -315 1725
rect -245 1725 -205 1735
rect -245 1715 -235 1725
rect -325 1705 -235 1715
rect -215 1715 -205 1725
rect -215 1705 -145 1715
rect -360 1695 -145 1705
rect -360 1670 -290 1675
rect -240 1670 -140 1675
rect -360 1665 -140 1670
rect -360 1660 -170 1665
rect -360 1655 -280 1660
rect -305 1650 -280 1655
rect -295 1645 -280 1650
rect -290 1640 -280 1645
rect -260 1655 -170 1660
rect -260 1645 -230 1655
rect -180 1645 -170 1655
rect -150 1645 -140 1665
rect -260 1640 -250 1645
rect -355 1625 -315 1635
rect -290 1630 -250 1640
rect -180 1635 -140 1645
rect -355 1605 -345 1625
rect -325 1605 -315 1625
rect -355 1595 -315 1605
rect -335 1575 -315 1595
rect -175 1575 -155 1635
rect -335 1565 -295 1575
rect -335 1495 -325 1565
rect -305 1495 -295 1565
rect -335 1485 -295 1495
rect -265 1565 -225 1575
rect -265 1495 -255 1565
rect -235 1495 -225 1565
rect -265 1485 -225 1495
rect -200 1565 -155 1575
rect -200 1495 -190 1565
rect -170 1495 -155 1565
rect -200 1485 -155 1495
rect -265 1450 -245 1485
rect -305 1440 -245 1450
rect -175 1445 -155 1485
rect -305 1430 -250 1440
rect -305 1405 -285 1430
rect -175 1425 -120 1445
rect -315 1395 -275 1405
rect -315 1225 -305 1395
rect -285 1225 -275 1395
rect -315 1215 -275 1225
rect -250 1395 -160 1405
rect -250 1225 -240 1395
rect -220 1225 -195 1395
rect -175 1225 -160 1395
rect -250 1215 -160 1225
rect -140 1270 -120 1425
rect -140 1185 -115 1270
rect -315 1090 -275 1100
rect -315 1030 -305 1090
rect -355 1020 -305 1030
rect -285 1020 -275 1090
rect -355 1010 -275 1020
rect -250 1090 -210 1100
rect -250 1020 -240 1090
rect -220 1030 -210 1090
rect -220 1020 -200 1030
rect -250 1010 -200 1020
rect -355 960 -335 1010
rect -375 940 -335 960
rect -310 960 -275 970
rect -310 920 -305 960
rect -375 900 -305 920
rect -335 895 -305 900
rect -310 890 -305 895
rect -285 890 -275 960
rect -310 880 -275 890
rect -250 960 -210 970
rect -250 890 -240 960
rect -220 920 -210 960
rect -220 900 -200 920
rect -220 890 -210 900
rect -250 880 -210 890
rect -235 790 -210 880
rect -235 785 -200 790
rect -315 775 -275 785
rect -315 715 -305 775
rect -355 705 -305 715
rect -285 705 -275 775
rect -355 695 -275 705
rect -250 775 -210 785
rect -250 705 -240 775
rect -220 715 -210 775
rect -220 705 -205 715
rect -250 695 -205 705
rect -355 280 -335 695
rect -315 645 -275 655
rect -315 585 -305 645
rect -310 575 -305 585
rect -285 575 -275 645
rect -310 565 -275 575
rect -250 645 -210 655
rect -250 575 -240 645
rect -220 575 -210 645
rect -250 565 -210 575
rect -295 460 -275 565
rect -240 535 -210 565
rect -235 520 -205 535
rect -225 510 -185 520
rect -225 490 -215 510
rect -195 490 -185 510
rect -225 480 -185 490
rect -295 440 -205 460
rect -290 400 -250 410
rect -290 330 -280 400
rect -260 330 -250 400
rect -290 320 -250 330
rect -275 280 -255 320
rect -365 270 -320 280
rect -365 200 -350 270
rect -330 200 -320 270
rect -365 190 -320 200
rect -295 270 -255 280
rect -295 200 -285 270
rect -265 200 -255 270
rect -295 190 -255 200
rect -225 280 -205 440
rect -225 270 -185 280
rect -225 200 -215 270
rect -195 200 -185 270
rect -225 190 -185 200
rect -365 180 -345 190
rect -400 160 -345 180
rect -365 130 -345 160
rect -205 170 -185 190
rect -205 160 -165 170
rect -205 140 -195 160
rect -175 140 -165 160
rect -380 120 -340 130
rect -270 125 -230 135
rect -205 130 -165 140
rect -270 120 -260 125
rect -380 100 -370 120
rect -350 110 -340 120
rect -290 110 -260 120
rect -350 105 -260 110
rect -240 105 -230 125
rect -350 100 -230 105
rect -380 95 -230 100
rect -380 90 -280 95
rect -400 60 -165 70
rect -400 50 -305 60
rect -315 40 -305 50
rect -285 50 -195 60
rect -285 40 -275 50
rect -315 30 -275 40
rect -205 40 -195 50
rect -175 40 -165 60
rect -205 30 -165 40
rect -380 20 -340 30
rect -380 0 -370 20
rect -350 0 -340 20
rect -380 -10 -340 0
rect -365 -35 -345 -10
rect -205 -35 -185 30
rect -365 -45 -320 -35
rect -365 -115 -350 -45
rect -330 -115 -320 -45
rect -365 -125 -320 -115
rect -295 -45 -250 -35
rect -295 -115 -285 -45
rect -265 -115 -250 -45
rect -295 -125 -250 -115
rect -225 -45 -185 -35
rect -225 -115 -215 -45
rect -195 -115 -185 -45
rect -225 -125 -185 -115
rect -280 -190 -260 -125
rect -415 -200 -320 -190
rect -415 -370 -400 -200
rect -380 -370 -350 -200
rect -330 -370 -320 -200
rect -415 -380 -320 -370
rect -295 -200 -250 -190
rect -295 -370 -285 -200
rect -265 -370 -250 -200
rect -295 -380 -250 -370
rect -280 -385 -260 -380
<< viali >>
rect -260 1940 -240 2010
rect -195 1225 -175 1395
rect -280 330 -260 400
rect -400 -370 -380 -200
<< metal1 >>
rect -360 2010 -110 2165
rect -360 1940 -260 2010
rect -240 1940 -110 2010
rect -360 1930 -110 1940
rect -360 1395 -110 1445
rect -360 1225 -195 1395
rect -175 1225 -110 1395
rect -360 1185 -110 1225
rect -325 790 -210 835
rect -325 785 -195 790
rect -375 400 -155 785
rect -375 330 -280 400
rect -260 330 -155 400
rect -375 315 -155 330
rect -355 280 -335 315
rect -225 280 -205 315
rect -425 -200 -70 -165
rect -425 -370 -400 -200
rect -380 -370 -70 -200
rect -425 -400 -70 -370
<< labels >>
rlabel locali -375 910 -375 910 7 D_bar
port 2 w
rlabel locali -375 950 -375 950 7 D
port 3 w
rlabel locali -360 1710 -360 1710 7 Q_bar
port 7 e
rlabel locali -360 1665 -360 1665 7 Q
port 6 e
rlabel metal1 -360 2040 -360 2045 7 GND
rlabel metal1 -425 -255 -425 -255 7 GND
port 1 w
<< end >>
