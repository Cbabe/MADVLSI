magic
tech sky130A
timestamp 1694559992
<< nwell >>
rect -130 165 270 315
<< nmos >>
rect -10 30 5 130
rect 185 30 200 130
<< pmos >>
rect -10 185 5 285
rect 185 185 200 285
<< ndiff >>
rect -60 115 -10 130
rect -60 45 -45 115
rect -25 45 -10 115
rect -60 30 -10 45
rect 5 115 55 130
rect 5 45 20 115
rect 40 45 55 115
rect 5 30 55 45
rect 135 115 185 130
rect 135 45 150 115
rect 170 45 185 115
rect 135 30 185 45
rect 200 115 250 130
rect 200 45 215 115
rect 235 45 250 115
rect 200 30 250 45
<< pdiff >>
rect -60 270 -10 285
rect -60 200 -45 270
rect -25 200 -10 270
rect -60 185 -10 200
rect 5 270 55 285
rect 5 200 20 270
rect 40 200 55 270
rect 5 185 55 200
rect 135 270 185 285
rect 135 200 150 270
rect 170 200 185 270
rect 135 185 185 200
rect 200 270 250 285
rect 200 200 215 270
rect 235 200 250 270
rect 200 185 250 200
<< ndiffc >>
rect -45 45 -25 115
rect 20 45 40 115
rect 150 45 170 115
rect 215 45 235 115
<< pdiffc >>
rect -45 200 -25 270
rect 20 200 40 270
rect 150 200 170 270
rect 215 200 235 270
<< psubdiff >>
rect -110 115 -60 130
rect -110 45 -95 115
rect -75 45 -60 115
rect -110 30 -60 45
<< nsubdiff >>
rect -110 270 -60 285
rect -110 200 -95 270
rect -75 200 -60 270
rect -110 185 -60 200
rect 85 270 135 285
rect 85 200 100 270
rect 120 200 135 270
rect 85 185 135 200
<< psubdiffcont >>
rect -95 45 -75 115
<< nsubdiffcont >>
rect -95 200 -75 270
rect 100 200 120 270
<< poly >>
rect -10 285 5 300
rect 185 285 200 300
rect -10 130 5 185
rect 185 130 200 185
rect -10 15 5 30
rect -35 5 5 15
rect -35 -15 -25 5
rect -5 -15 5 5
rect -35 -25 5 -15
rect 185 15 200 30
rect 185 5 225 15
rect 185 -15 195 5
rect 215 -15 225 5
rect 185 -25 225 -15
<< polycont >>
rect -25 -15 -5 5
rect 195 -15 215 5
<< locali >>
rect -105 270 -15 280
rect -105 200 -95 270
rect -75 200 -45 270
rect -25 200 -15 270
rect -105 190 -15 200
rect 10 270 50 280
rect 10 200 20 270
rect 40 200 50 270
rect 10 190 50 200
rect 90 270 180 280
rect 90 200 100 270
rect 120 200 150 270
rect 170 200 180 270
rect 90 190 180 200
rect 205 270 245 280
rect 205 200 215 270
rect 235 200 245 270
rect 205 190 245 200
rect 30 170 50 190
rect 220 170 240 190
rect 30 150 250 170
rect 220 125 240 150
rect -105 115 -15 125
rect -105 45 -95 115
rect -75 45 -45 115
rect -25 45 -15 115
rect -105 35 -15 45
rect 10 115 50 125
rect 10 45 20 115
rect 40 45 50 115
rect 10 35 50 45
rect 140 115 180 125
rect 140 45 150 115
rect 170 45 180 115
rect 140 35 180 45
rect 205 115 245 125
rect 205 45 215 115
rect 235 45 245 115
rect 205 35 245 45
rect 25 15 45 35
rect 140 15 160 35
rect -115 5 5 15
rect -115 -5 -25 5
rect -35 -15 -25 -5
rect -5 -15 5 5
rect 25 -5 160 15
rect 185 5 225 15
rect -35 -25 5 -15
rect 185 -15 195 5
rect 215 -15 225 5
rect 185 -25 225 -15
rect 185 -45 205 -25
rect -115 -65 205 -45
<< viali >>
rect -95 200 -75 270
rect -45 200 -25 270
rect 100 200 120 270
rect 150 200 170 270
rect -95 45 -75 115
rect -45 45 -25 115
<< metal1 >>
rect -115 270 255 280
rect -115 200 -95 270
rect -75 200 -45 270
rect -25 200 100 270
rect 120 200 150 270
rect 170 200 255 270
rect -115 190 255 200
rect -115 115 255 125
rect -115 45 -95 115
rect -75 45 -45 115
rect -25 45 255 115
rect -115 35 255 45
<< labels >>
rlabel metal1 -115 80 -115 80 7 VN
port 5 w
rlabel locali -115 -55 -115 -55 7 B
port 2 w
rlabel locali -115 5 -115 5 7 A
port 1 w
rlabel locali 250 160 250 160 3 Y
port 3 e
rlabel metal1 -115 240 -115 240 7 VP
port 4 w
<< end >>
